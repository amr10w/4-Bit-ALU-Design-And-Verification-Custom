module simple_print;
  
endmodule
